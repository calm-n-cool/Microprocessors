`timescale 1ns / 1ps

module BUS(input [7:0] in,output [7:0] out);
assign out = in;
endmodule
